`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.12.2022 11:25:34
// Design Name: 
// Module Name: NN_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module NN_tb;
    
    logic signed [7:0] test_data_b [0:783] = '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 116, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 90, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 76, 105, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 127, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 127, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 122, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 99, 127, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 127, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 115, 127, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 127, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 127, 108, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 127, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 43, 89, 124, 127, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 127, 42, 0, 0, 0, 23, 24, 58, 72, 75, 120, 121, 117, 89, 120, 126, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 126, 118, 103, 103, 103, 126, 127, 125, 120, 99, 71, 45, 14, 2, 116, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 88, 88, 88, 88, 88, 49, 28, 0, 0, 0, 0, 0, 51, 127, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 127, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 127, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 127, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 127, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 127, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 127, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 127, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 127, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 };
    logic signed [7:0] test_data_a [0:783] = '{ 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 40, 103, 127, 127, 127, 127, 48, 40, 40, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 79, 79, 79, 84, 126, 126, 126, 126, 126, 126, 126, 126, 126, 105, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 120, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 126, 126, 126, 119, 56, 107, 126, 126, 126, 126, 126, 126, 126, 126, 126, 105, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 17, 17, 17, 15, 0, 15, 74, 17, 102, 117, 126, 126, 126, 126, 126, 118, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 17, 99, 126, 126, 126, 126, 122, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 16, 101, 101, 108, 126, 126, 126, 126, 120, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 83, 126, 126, 126, 126, 126, 126, 126, 119, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 126, 126, 126, 126, 126, 126, 126, 126, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 100, 126, 126, 126, 126, 126, 126, 126, 115, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 43, 43, 43, 124, 126, 126, 126, 126, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 76, 126, 126, 126, 125, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 119, 126, 126, 126, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 116, 126, 126, 75, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 101, 126, 126, 126, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 105, 105, 105, 29, 18, 18, 10, 13, 18, 75, 111, 126, 126, 126, 126, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 126, 126, 126, 126, 126, 126, 97, 107, 126, 126, 126, 126, 126, 126, 78, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 118, 117, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 78, 123, 126, 126, 126, 126, 126, 126, 126, 126, 79, 78, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 126, 126, 126, 126, 126, 63, 39, 39, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 };
    
localparam period = 20;

reg clk, enable, reset;  
reg signed [7:0] img [0:783];
reg [7:0] digit_out;
reg NN_done;

    neural_network NN(.clk(clk), .enable(enable), .reset(reset)
                  .img(img), .digit_out(digit_out), .NN_done(NN_done));

initial begin
clk = 0;
enable = 0;
reset = 0;
img = test_data_a;
#145
enable = 1;
end

always begin
#10 clk = ~clk;
end

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.12.2022 22:18:50
// Design Name: 
// Module Name: avg_pooling
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


/**********
* Average pooling implementation
*
* Inputs: clk => clock signal, pool_en => enable signal, 
*         in1 => top left pixel value, 
*         in2 => top right pixel value,
*         in3 => bottom left pixel value,
*         in4 => bottom right pixel value,
*
* Outputs: out => in pixels average
*          pool_done => done signal
* 
***********/

module avg_pooling(
    input clk,
    input pool_en,
    input [7:0] in1,
    input [7:0] in2,
    input [7:0] in3,
    input [7:0] in4,
    output [7:0] out,
    output  pool_done
    );
    
    reg [15:0] pool_out;
    
    always @(posedge clk) begin
        if(pool_en == 1) begin
            pool_out <= (in1+in2+in3+in4)>> 2; //Calculate average
        end
        
    end
    
    assign out = pool_out[7:0];
    assign pool_done = (pool_out==(in1+in2+in3+in4)>> 2)? 1:0;

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.01.2023 23:47:02
// Design Name: 
// Module Name: dense_layer
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/**********
* Dense layer implementation
*
* Parameters: NEURON_NB => The # of neurons
*             IN_SIZE => The input vector size
*             WIDTH => The width of the weights and biases
*
* Inputs: clk => clock signal, layer_en => enable signal, 
*         reset => active high sync reset signal, in_data => in vector, 
*         weights => neurons weights, biases => neurons biases
*
* Outputs: neuron_out => dense layer output
*          layer_done => done signal
* 
***********/

module dense_layer # (parameter NEURON_NB=32, IN_SIZE=196, WIDTH=8)(
    input clk,
    input layer_en,
    input reset,
    input signed[2*WIDTH-1:0] in_data [0:IN_SIZE-1],
    input signed[WIDTH-1:0] weights [0:NEURON_NB-1][0:IN_SIZE-1],
    input signed[WIDTH-1:0] biases [0:NEURON_NB-1],
    output signed[4*WIDTH-1:0] neuron_out [0:NEURON_NB-1],
    output layer_done
    );
    
    reg [0:NEURON_NB-1] neuron_done;
    reg done = 0;
    
    neuron #(.IN_SIZE(IN_SIZE), .WIDTH(WIDTH)) dense_neuron[0:NEURON_NB-1] (.clk(clk), .en(layer_en), .reset(reset), 
                                                                            .in_data(in_data), .weight(weights), .bias(biases), 
                                                                            .neuron_out(neuron_out), .neuron_done(neuron_done)); // Neuron submodules
    always @(posedge clk) begin
        if(neuron_done == '1) begin //All neurons done
            done <= 1;
        end
    end
    
    assign layer_done = done;

    
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.12.2022 09:16:01
// Design Name: 
// Module Name: dense_layer1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/**********
* 1st dense layer implementation (hidden layer)
*
* Inputs: clk => clock signal, enable => enable signal, 
*         reset => active high sync reset, pooled_img => in vector, 
*
* Outputs: layer_out => dense layer output
*          layer_done => done signal
* 
***********/


module dense_layer1(
    input clk,
    input enable,
    input reset,
    input signed [15:0] pooled_img [0:195],
    output signed [15:0] layer_out [0:31],
    output layer_done
    );
    
    reg signed [31:0] dense1_res [0:31];
    reg signed [15:0] relu_res [0:31];
    
    //Biases and weights
    localparam signed [7:0] B_ARRAY_L2 [0:31] = '{ 21, -2, -5, 6, 12, -16, 6, 1, 17, 8, 3, 5, -23, 17, 8, 5, 5, 22, 8, 8, 1, 6, -9, 9, 15, 20, -13, -5, 2, 7, 12, 24 };
    
    localparam signed [7:0] W_ARRAY_L2 [0:31] [0:195] = '{
    { 7, -1, 9, 12, 17, 36, 29, 35, 33, 44, 25, 23, -8, 7, 0, 11, -10, -4, -6, 5, 5, 28, 27, 29, 12, 28, 1, 9, -1, -11, -41, -26, -8, -22, -22, 6, -1, 12, 16, 14, -11, 12, -8, -31, -31, -2, -21, -7, 11, 5, 1, -2, -26, 1, 4, -14, -5, -4, -44, -20, -2, 6, 20, 10, -3, -31, -26, -28, -5, -18, -3, -15, -44, 1, -1, -12, 1, 14, -16, -17, -1, 2, 28, -28, 7, 2, -16, 9, -7, -8, -1, -5, -4, 7, 10, 12, 25, -41, 10, 4, 4, -2, 0, 8, 6, -12, -26, -7, 3, 7, 31, -18, -11, 9, 6, -19, 9, 29, 6, -9, -17, -18, -1, -3, 24, -25, 15, -7, -15, -12, 14, 12, -5, -6, 5, -7, 4, 5, 23, -25, 3, 0, 6, -1, 21, 32, 13, 14, 17, 10, 5, 13, -8, 11, 2, -1, 10, 18, 10, 16, 14, 14, 11, 1, -20, -23, -24, 20, 0, -28, -2, -13, -9, 1, -16, -29, -32, -17, -37, -43, -6, 18, -1, -1, -29, -39, -56, -33, -52, -46, -56, -41, -33, -16, -5, 1 },
    { -6, -9, 2, -6, 2, -15, -22, 8, -20, 23, 25, 17, -9, 4, -2, 9, 18, 17, -18, -6, -23, -8, 8, 27, 33, -1, -11, -9, -5, 12, 21, 1, -12, -4, 3, 14, 14, 6, -4, -5, -10, 1, 25, 9, 23, -3, -6, -17, 5, 24, 12, -10, -18, -5, 9, 27, -17, 1, 5, -8, -16, -45, -9, 30, -7, -23, -18, -33, 6, 18, -11, -20, -36, -29, -26, -2, 45, 32, -4, -15, -37, -56, -27, 4, -20, -28, -22, -10, 27, 33, 29, -29, -14, -19, -6, -5, -62, -29, -8, -15, -16, 1, -11, -3, -14, -20, 2, 10, 22, 27, -20, -50, 11, -3, 13, 7, -1, 1, 2, -8, 2, 3, 11, 31, -19, -55, -16, 16, 8, 13, 5, 7, 17, 13, 6, 6, -9, 8, -6, -28, 4, -6, -10, 0, 0, -8, -1, 7, 3, 10, -16, -4, 9, -15, 20, 1, -15, -16, -11, 12, 3, -7, -1, 0, -9, -5, -12, 27, 5, 8, 16, 33, 33, 3, -6, -2, -3, 19, 12, 11, 22, 20, 4, -4, 7, -12, -34, -42, -56, -12, 17, 0, 0, -13, 8, -7 },
    { 8, 8, 1, -8, 5, -2, -16, 14, -10, -13, -14, -5, 2, 8, 4, 12, -18, 9, -6, 4, 15, 1, -1, -17, -30, -6, -3, -20, 6, 28, 21, 12, 1, 17, 8, 9, -6, -13, -8, -14, -12, 2, -27, 9, -15, -8, 1, -9, -1, 4, 5, -26, -14, -23, -4, -10, -40, 5, 22, 3, -5, -19, 5, 23, 27, -1, -31, -38, -29, 21, -18, 12, 18, 15, 0, 24, 13, 34, 36, 20, -46, -49, -29, 12, -26, -2, 10, -3, 9, 3, 12, 39, 46, 2, -47, -40, -5, 2, -16, 5, -28, -25, -23, -17, 7, 29, 21, -32, -42, -26, 1, 40, 16, -6, -41, -35, 3, -11, 9, 7, -22, -39, -15, -14, 7, 40, -27, -8, -37, -21, -2, -4, -4, -4, -6, 1, 10, -3, -13, 18, 10, -10, -22, 2, 3, -7, -16, 5, 8, 21, 6, -2, 13, 17, 14, 25, -10, 0, -7, -2, -3, 2, -3, 12, 13, 11, 15, 3, 8, -17, -16, -20, -10, -11, -5, -1, 5, 16, 17, -8, 8, 25, 1, 15, -19, 0, 8, -9, -15, -3, -1, 3, -11, -23, -3, -6 },
    { 2, -1, -8, -23, -29, -47, -51, -28, -3, -28, -34, -32, 7, -7, -5, -12, 11, -2, -25, -25, -47, -62, -45, -38, -31, -8, 18, 11, -5, 23, 41, 14, 17, 4, 1, -9, -21, -16, -16, 8, 9, -2, 29, 31, 23, 21, 33, 45, 30, -14, -16, -9, -1, 12, -9, 1, 29, 6, 8, 10, 21, 30, 22, -4, -5, 6, 8, 14, -49, -5, 0, -4, -20, -27, -24, -25, -21, -11, 3, 6, 10, -1, -41, -22, 15, -20, -49, -45, -33, 2, -11, -13, 1, -4, -6, -23, 11, 13, -2, -32, -19, -4, -5, 17, -5, 0, 10, 19, 10, 9, 20, 54, 2, -26, -23, 5, 20, -19, 7, 10, 4, 25, 12, 4, 26, 54, 19, 6, -2, 0, -15, -4, 19, 4, 0, -7, -7, 3, 2, 35, 9, 24, -4, -11, -4, 10, 5, 7, -20, -44, -18, -1, -15, 20, 2, -1, -6, 7, 0, 5, 10, 4, -4, -23, -10, -5, -15, -6, -6, 6, 7, 11, -8, 7, 2, 6, -8, -35, -46, -20, 5, 1, -9, -19, -28, -8, 5, 0, -15, 3, 21, -7, -26, 11, -1, 5 },
    { -9, 4, 3, 4, 2, 2, 3, -3, 9, 10, 13, 8, 9, 2, 4, 9, -25, -31, -21, -33, -24, -14, -30, -9, -18, 15, 13, -1, 0, 5, -30, -27, -31, -14, -11, -8, -7, -4, -3, -11, 11, 7, -7, 3, -3, -5, -3, -5, 1, 9, 7, 18, 19, 12, 9, -7, 24, 7, 15, 2, 6, 20, 24, 21, 19, 19, 20, 31, 19, 26, 25, 7, 19, 25, 23, 27, 36, 9, 1, -5, -9, 6, 32, 64, 35, -2, 4, -5, 3, -17, -26, -32, -18, -16, -15, -18, 13, 30, 16, -25, -37, -33, -30, -26, -20, -20, -11, -12, -14, -1, -1, 24, -12, -3, -19, -18, 2, 3, 9, -9, -3, -31, -16, -28, -1, 39, 21, -16, -4, 13, 18, 3, 3, 1, -5, -7, -17, -13, -3, 27, -6, -5, 0, 8, 8, 0, 4, 8, 5, 19, 9, 7, 30, 27, -13, -25, 11, -4, -3, -2, 10, 9, 10, 7, -3, 19, 33, -23, 6, 0, -12, -20, 5, 3, 22, 38, 37, 43, 11, 14, 36, 3, 0, -6, -20, -18, 23, 20, 26, 39, 32, 42, 14, 14, -3, -2 },
    { -8, -1, 6, 18, 35, 26, 34, -13, 12, 43, 26, 22, 9, 0, -8, -11, 10, 32, 46, 35, 38, 17, -2, -3, 7, -4, -26, 2, -1, -5, 12, 6, -3, -14, -17, -23, -15, -4, -13, -17, -15, 32, 31, 8, -16, -4, 7, -2, 4, 18, 6, -4, -6, -8, 17, 0, 1, 3, 6, 15, 21, 17, 13, 5, -14, -8, 16, 12, -9, 20, -16, 35, 12, 20, 9, -17, -40, -30, -5, 28, 31, 23, -29, -34, -2, 18, 10, -13, -25, -30, -21, 13, 35, 21, 19, 27, 7, -54, -2, -4, -13, -8, -13, 2, 17, 29, 4, 11, 8, 0, 3, -36, 33, 24, 9, 5, -8, 8, 23, 10, 12, 0, -11, -3, 8, -18, 6, 16, 16, -6, -22, -1, 8, 8, 14, 5, -14, -24, -33, 0, -5, -14, -7, 12, 0, -15, -4, 19, -4, -5, -23, -30, -16, -12, -6, 7, -2, -8, -15, -2, -16, -15, -9, -16, -21, -4, -19, -21, -2, 24, 23, 24, 18, 15, 0, 10, 1, 4, 12, 0, -2, -10, -7, 17, 25, 69, 72, 49, 45, 45, 36, 33, 35, 44, -4, 2 },
    { 7, -9, -9, -6, -8, -13, -37, -17, -32, -17, -11, 8, 9, 7, -4, -2, -1, 5, 21, 10, 4, -12, -19, -3, 17, 1, 17, 11, 9, 29, 26, 22, 5, 11, 7, 9, -1, 1, -2, 10, 26, 41, 35, 13, 13, -5, 9, 9, 7, -5, 10, 9, 5, 1, 39, 47, 17, 10, 13, 17, 12, 16, 30, 27, 2, 4, 4, 10, 6, 12, 34, 13, 22, 8, 6, 12, 14, 5, -16, -16, -34, -36, -41, 27, 23, -10, 0, -13, -11, -11, -29, -9, 4, 7, -25, -55, -72, 20, 29, 11, -29, -32, -28, -43, -29, 1, -2, 14, -5, -1, 4, 49, 9, 9, -35, -38, -29, -42, -21, -2, 0, 15, 12, 13, 38, 66, 27, 34, -12, -6, 2, -34, -1, 19, 11, 2, 9, 10, 27, 56, -10, 29, -4, 7, 5, 19, 28, 19, 12, 2, -2, 7, 9, 17, 11, -4, 16, 13, 10, 15, 2, 8, 9, -4, -8, -12, -2, 25, -6, 17, 33, 16, 18, 4, 11, -1, -8, 6, -16, -33, -26, 16, -5, -7, -23, 11, 13, 3, 12, 23, 26, 32, 4, -9, -3, -5 },
    { -4, -5, -2, -20, -24, -6, 1, -8, 7, -45, -31, -26, 8, 1, 4, 12, -8, -4, -22, -4, 3, -2, -7, -21, -17, -17, -3, -4, 9, 9, 27, 24, 25, 5, 6, 10, 18, 22, 4, 2, -9, -15, 36, 52, 46, 21, -11, 3, 12, -6, -1, 15, -6, 23, 0, -1, 27, 75, 36, 1, -2, 10, 18, 6, 15, 34, 24, 25, -6, -11, 33, 44, -9, -20, -3, -7, 8, -22, 7, 14, 23, 14, -29, -56, 26, 12, -19, 0, 5, 14, 3, -29, -23, -5, -22, 1, 11, -29, 7, -14, 5, 9, 13, 3, -15, -17, -7, 29, 15, 18, 21, 16, 26, -15, 1, 2, 15, -6, 3, -9, 11, 12, 13, 27, -5, 10, 20, 9, 12, -3, 3, -6, -6, -5, 11, 3, 10, 4, -22, -8, 26, 12, 5, 2, 6, 9, 14, 2, -13, -12, -20, -24, -60, 10, -3, 1, -21, 22, 9, 15, 19, 12, 6, 2, -12, -28, -26, -19, -8, 32, 10, 17, 5, 4, 11, 7, -9, -33, -46, -35, -14, -17, -8, -5, -19, -5, -20, -26, -29, -43, -14, -8, -34, -5, 3, -9 },
    { -2, 1, 0, -23, -20, -37, -24, -20, -42, -34, -34, -15, -2, -1, 7, -14, -9, -44, -38, -29, -16, 6, 18, 7, -16, -45, -29, -17, 1, 25, -16, -21, -1, 3, -11, -1, 20, 24, 14, 1, -21, -17, 23, 10, -23, -17, -18, -19, -32, -27, 7, 23, 8, 15, -13, -7, -28, 13, -24, -29, -20, -4, -9, -49, 17, 27, 16, 15, -12, 5, -13, -6, -25, -17, -11, -8, -23, -41, 27, 30, 0, -29, -14, 28, -12, -11, -12, -18, -18, -25, -15, -8, 8, 19, -5, -32, -3, 46, 4, 24, 20, 23, 15, 3, 3, -13, 13, -2, -11, -16, 10, 50, 32, 39, 41, 22, 18, 22, 30, 4, 14, 1, 1, -9, -5, 42, -4, 46, 35, 27, 11, 19, 12, -3, 2, 11, -9, -17, 5, 8, -23, 37, 9, 0, -13, -14, -23, -7, 21, 14, 6, 12, 18, -14, 5, 26, 20, -13, -16, -19, -21, -5, -7, 17, 34, 15, 22, -2, -4, -4, -19, -5, -12, -10, 1, 8, 7, 5, 16, 18, -17, 19, -3, 4, 17, -1, 2, 7, 24, -14, -33, -41, 5, 5, -10, -1 },
    { 6, 7, 13, 12, 21, 8, 3, 1, 31, 28, 25, 26, 1, 0, 3, 7, 5, 16, 26, 26, 11, 12, 11, 5, -9, 23, 0, 12, 2, -5, -8, -6, 1, 18, 23, 15, 13, 10, -1, -18, -20, 7, -36, -22, -8, -17, 3, 19, 24, 21, -2, -11, -7, -5, 2, -18, -26, -16, -4, -12, -10, 8, -6, 0, -21, -14, 3, -7, -19, -3, -43, -28, 10, 2, 8, 0, -4, -7, -23, -3, 13, 15, 19, -19, -28, -4, 13, 1, 2, -10, 0, -10, -6, 2, 28, 23, 9, 9, -24, 4, -10, 1, -1, 14, 15, 12, 11, 7, 5, -11, -9, 28, -17, 6, 0, 11, 12, 17, 25, 23, 8, 7, -13, -1, 8, 29, -19, -6, 7, 28, 21, 19, 20, 17, 21, 7, -8, 11, 6, 5, -7, 20, 16, 16, 20, 16, 12, 16, 20, 9, 7, 12, 16, 2, -13, 22, -6, -12, -1, 4, 12, 3, 0, 4, 14, 37, 16, -26, 1, -36, -44, -25, -17, -11, -8, -8, -5, 7, 10, 13, 28, 7, -1, 10, 33, 21, 12, 16, 21, 13, 5, 0, 1, -9, 19, 2 },
    { 6, 3, 3, -2, -7, 13, 7, 11, -3, 42, 36, 26, -5, 5, -5, 9, 23, 14, -8, -44, -47, -19, -6, 6, 10, 34, 4, -1, 7, 3, -2, -41, -25, -30, -15, -8, -3, 3, 5, 2, -8, 22, -30, -11, -8, -19, -34, -17, -14, 1, 2, 13, 14, 11, -2, -9, -33, -27, -13, -21, -36, -13, 12, 11, -6, -7, 4, 17, 9, -5, 1, -41, -2, -48, -34, 17, 39, 17, -14, -14, 2, 6, -13, -4, -10, -25, -11, -20, -19, 3, 24, 24, 19, -10, 17, 25, -26, -41, -10, -21, -42, -22, -5, -1, 8, 25, -1, -11, -16, -30, -38, -49, -11, -28, -28, -5, 22, 11, 14, 5, -19, -18, 2, -18, -21, -31, -9, -51, -28, -10, 17, 16, 6, -21, -16, -10, 10, -22, -11, 10, 14, -59, -20, -6, 1, 7, -1, -20, -22, 0, -1, -18, -9, -7, 2, -22, -10, 0, -7, 3, 17, 11, 2, -3, -15, -19, 14, 12, -6, -39, -28, -8, -2, -1, 1, 6, -1, -2, 1, -24, -7, -7, 6, 18, 13, 8, 6, 0, 13, 18, 31, 5, 19, -14, 5, 3 },
    { 8, 1, 6, 9, -8, 15, 8, -8, 32, 21, -10, -6, -5, 8, -1, -11, -3, 46, 38, 51, 52, 33, 6, -10, -14, 5, 23, 1, 10, 13, 10, 10, 9, 13, -1, 10, 5, 1, -14, -14, -23, 7, 35, 26, 18, 1, 9, 15, 10, 17, 6, 11, -2, -1, -40, -13, 21, 34, 0, -4, -8, -32, -51, 5, 32, 7, 0, -2, -64, -38, 10, -5, -34, -61, -81, -56, -50, -2, 7, 6, -1, 2, -30, -20, -8, -16, -44, -35, 5, 20, 15, -1, -13, -11, 10, 6, -20, -10, -11, -2, 17, 28, 31, 18, 4, -8, -11, -17, 7, -2, -18, 35, 12, 20, 14, -4, 2, 3, -2, -9, 2, 6, -9, -12, -15, 43, 27, 8, -16, -11, 0, -10, 11, 3, 12, -4, -5, -17, -11, 24, 10, 27, -4, -6, -7, 7, 26, 20, 9, 9, 5, 12, 12, 50, 13, 41, 2, 7, 11, 18, 5, 12, -4, 4, 5, 16, 24, 22, 7, 20, 5, 7, 13, 12, 21, -1, 1, -10, -13, 6, 25, -3, -3, 5, 5, -3, -8, 22, 18, 4, -4, 5, -16, -3, 7, -8 },
    { -7, 3, 4, 14, 24, 25, 20, -6, 25, 42, 27, 12, -2, 8, 5, 15, 15, 16, 41, 40, 34, 10, 9, 24, 27, 4, 2, -21, 7, 9, -2, 8, 1, 11, 1, 21, 27, 22, 24, -22, 3, 38, 18, 6, 9, 6, -2, -4, 11, 15, 14, 11, -1, -4, -4, -9, -19, 12, 5, -2, -5, -7, 9, 14, 0, 12, 21, 16, 1, 8, -27, 9, 0, -5, -20, -6, 31, 22, 0, 17, 10, 12, 21, 15, -30, -6, 8, -17, -24, 0, 38, 26, 16, 8, -7, -9, 6, 14, 4, -19, -22, -17, -9, 16, 23, 1, 3, 8, -10, -24, -1, -15, 15, 4, 1, -12, 7, 21, -6, -24, 13, 5, -14, 0, -7, -20, -9, 1, 16, 22, 29, 11, -15, -1, 6, 1, -2, 8, -52, -37, 20, -3, 2, 21, 6, 4, 12, 13, 9, 2, 13, -6, -50, -19, -1, 19, -20, -11, -1, 11, 26, 16, 19, 4, -6, 7, -30, -38, -8, 11, -23, -7, 9, 23, 24, 24, 16, 2, -1, 0, -9, -13, -1, -3, 10, 17, 4, 18, 17, 11, 8, 12, -2, -11, 10, -2 },
    { 3, 5, 1, 2, 0, 14, 20, 0, -12, -11, -3, -12, 1, 7, -4, 5, -10, -8, -50, -33, -10, -9, -10, -13, -7, 10, -20, -10, 1, -11, -13, -25, -38, -7, 9, 5, -4, -5, -4, 6, 16, -1, -38, -25, -5, -33, -10, 13, 6, 0, -18, 0, -5, 4, 34, 38, -21, -40, -45, -24, -4, 1, 1, -10, -13, 1, 13, 11, 58, 24, -10, -31, -55, -40, -3, 9, 12, 3, -8, -10, 2, 17, 46, 18, -5, -25, -48, -27, 2, 28, 41, 25, 12, -19, -17, -12, -20, -20, 6, -6, -28, -34, 2, 22, 26, 25, 14, -7, -11, -27, -32, -45, 4, -7, -8, -17, -25, -14, 15, 22, 14, -15, -27, -38, -26, -33, -29, -17, -3, -15, -22, -31, -1, 20, 10, -6, -23, -39, -23, 21, -5, -16, -10, -8, -8, -7, -3, 9, 9, -8, -41, -46, -38, 0, -8, -15, 18, -5, 9, 8, 20, 5, -2, -34, -47, -31, -10, 10, -7, -17, -7, -9, 15, 22, 19, 0, -11, -15, -13, 19, 13, 2, 7, 5, -13, -36, -35, -14, -21, -17, -7, -8, -3, 11, 1, -1 },
    { 3, 8, -8, -19, -28, -35, -22, -38, -31, -38, -24, -28, -1, -1, -3, -15, -30, -60, -60, -71, -127, -106, -80, -53, -35, -23, -28, -12, 2, 12, 0, -1, -32, -20, -9, -10, -14, -21, -14, 7, 13, -25, -21, 35, -17, -1, 15, 14, 9, 16, 6, 6, 8, 2, -3, 14, -3, 8, 9, 22, 14, 1, 0, 6, -1, 3, 7, 0, -4, 6, -6, 18, 23, 22, 18, 17, 12, 6, 13, 10, 24, -6, -27, -3, 15, 26, 9, 5, 15, 16, -20, 13, 22, 15, 35, 0, -20, 3, 0, 37, -3, 5, 7, -6, -15, 18, 27, 21, 21, 4, -29, 4, -16, 1, -19, 3, 1, -8, 7, 15, 17, -4, -6, -11, -33, 4, 8, -6, -37, -20, -15, -20, 1, -3, -18, -33, -19, -51, -49, 8, -15, -45, -25, -28, -7, -13, -4, -10, -10, -18, -30, -26, -8, -28, 0, -27, -28, 3, 0, 2, 4, -6, -10, -7, 6, 1, -7, -29, -2, 1, 20, 20, 7, 2, -13, -9, -15, -11, 21, 9, -13, -7, -3, 18, 26, 44, 45, 9, 13, 33, 18, 12, 4, 10, 18, 0 },
    { 8, -2, -8, -18, -29, -16, -3, -13, -17, -34, -34, -32, 5, -5, 5, -2, -11, -46, -44, -32, -31, -11, -10, -17, -23, -33, -2, 11, 3, -32, -5, -28, -34, -3, 9, 6, -4, -15, -18, -42, -8, 23, -22, 23, -34, -25, -8, 13, 17, 15, 25, 14, 8, -9, -13, -2, 4, 8, -23, 3, 1, 6, 15, 19, 9, 24, 18, 10, 20, 23, 20, 9, 6, 6, 14, 11, 18, 15, 13, 21, 23, 28, 0, 7, 16, 28, 31, 17, 13, 7, -9, -8, 0, 23, 28, 14, -21, -3, 10, 11, 5, 19, 11, 8, -5, -22, 6, 25, 9, -5, -18, -13, -14, -20, 1, 6, 4, 2, 0, 1, 21, 1, -1, -12, -22, -19, 28, -17, -11, -6, -15, -3, -16, 7, 5, -1, -11, -28, -24, -5, 14, -26, 13, -5, -16, -13, -14, -21, -9, -21, -24, -30, -3, -22, -16, -1, -15, 14, 7, 12, -4, -9, -24, -37, -27, -3, -3, -19, 4, 32, 26, 20, 11, 13, 7, 3, -7, 3, 6, -2, -14, -19, 8, 17, 14, 43, 64, 41, 49, 45, 41, 29, 33, 26, 13, 4 },
    { 1, 3, -3, -12, 24, -5, 8, 18, 11, 11, 4, -14, 5, 9, -3, -5, 22, 21, 3, -8, 28, 47, 38, 35, 36, -2, 2, 13, -4, 3, 9, 16, 8, 10, -2, 2, -5, -1, 18, 24, 17, 7, 2, -5, 3, 4, 3, 8, 9, 10, 2, 8, 13, -1, 42, 5, 32, 4, -11, 3, 2, 12, 31, 0, -7, -8, -11, -8, 18, -7, 55, 12, -5, -2, 5, 26, 13, -20, 6, -13, -19, -20, -17, -5, 34, 9, 21, 17, 9, -1, -40, -16, 7, -1, 4, 18, -30, -35, 24, 12, 29, 19, 22, -10, -27, -14, 0, 3, 19, 22, -4, -31, 13, -3, 0, 5, 21, 3, -28, -5, -7, 14, 7, 4, -13, -34, 14, 2, -10, -10, 7, -10, -66, 18, 20, 22, 19, -1, -4, -36, -17, -3, -2, -9, 2, -14, -16, 33, 41, 18, 15, -5, 19, -15, 3, -14, -5, -18, -19, -18, 1, 32, 23, 15, 4, -13, 14, 13, -1, 26, 9, -16, -24, 3, 4, 9, 21, 13, 10, 7, -3, -20, 3, -1, -14, 15, 56, 33, 37, 59, 79, 73, 94, 52, 16, -1 },
    { 6, -8, -4, -5, -12, 11, 0, 3, 13, -32, -37, -26, 6, -2, -4, 10, -13, -24, -16, -14, 2, 0, 15, 2, -8, -14, -1, -5, -12, -19, -57, -27, -12, 5, 6, 21, 17, 9, 12, 4, 1, 5, -36, -35, -23, 6, 1, 22, 3, 5, 12, 10, 6, 20, 8, -11, 2, -16, -17, -1, 19, 16, 3, 4, 14, 1, 12, 19, 53, -11, 2, -7, 10, 18, 16, 9, 6, 3, -5, 14, 17, 24, 33, 10, -10, 8, 9, 26, -1, 7, 0, -29, -6, 5, 11, 16, 17, -8, -5, -22, 7, 13, 15, 6, -8, -41, -20, -12, 0, 12, 13, -33, -23, -1, 7, 6, 13, 0, -22, -19, 4, -6, -8, 5, -8, -14, 8, -9, 17, 24, 11, 16, 6, 2, -7, -4, -3, 2, 6, -33, 3, 14, 10, 14, 16, 11, 16, -1, 2, -9, 10, 7, -15, 18, -6, -16, 1, 10, 16, 14, 11, 12, 2, 2, -4, 2, -13, 10, -5, -9, -18, -29, -3, 0, 1, 12, 10, 12, -5, 15, 9, -7, -8, 6, -40, -53, -49, -35, -13, -14, -18, -2, -3, 2, -9, -1 },
    { 2, 6, -11, -21, -14, -32, -42, -21, -17, -21, -30, -17, -8, 7, -7, -3, -21, -25, -56, -76, -57, -45, -23, 5, -7, -7, -9, -19, -3, 1, -1, 2, -17, -1, -12, -11, 1, -4, 5, 14, 5, 11, 9, -18, 22, 16, 27, 7, -13, -8, -3, -6, -15, 5, 11, 13, -39, 3, 11, 25, 22, 10, 9, -8, 13, -3, 8, 20, 55, 45, -37, -8, 14, 11, 26, 16, -9, -25, -9, -7, -4, 19, 41, 61, -20, -22, 11, 20, 18, 34, 21, -3, -13, -5, 16, -2, 0, 44, 12, -12, -2, 4, 28, 45, 46, 30, 18, 0, -5, -5, -3, 28, 4, 7, -32, -21, -8, 5, 32, 33, 10, -8, -8, 14, -1, 9, -18, -4, -9, -28, -47, -35, -33, -15, -3, -20, 0, 2, 0, -19, -2, 11, 1, -11, -17, -24, -31, -12, -3, -3, 8, 23, 6, -13, -8, 28, 2, 2, 1, 12, -2, -7, -4, 8, 11, 18, 5, 21, 3, 23, -7, 10, 25, 37, 26, 28, 18, 15, 11, 12, 7, -22, 1, -14, -13, -32, -37, -11, -5, -19, -11, -21, -13, -11, -19, 1 },
    { 3, 7, 9, 12, 21, 9, 13, -6, 40, 31, 32, 23, 1, -6, 3, 5, 33, 31, 29, 27, 17, 19, 26, 38, 50, 21, 14, 7, 6, 11, -1, 3, 8, -3, -9, 6, 7, 0, 6, 7, 13, 36, 24, 18, 21, 8, -12, -32, -36, -30, -30, -35, -36, -25, 30, 5, 42, 25, 13, 1, -2, -18, -27, -38, -22, -23, -5, 1, 8, 3, 32, 24, 13, 2, 12, 30, 28, 20, 11, 6, 12, -1, 24, 8, 14, 32, -10, 10, 27, 25, 13, 19, 11, 9, -6, 11, 27, 0, 17, 19, 0, 10, 7, 3, 1, 5, 11, 20, 12, 36, 28, -40, 16, 20, 16, -2, -14, -4, -1, 7, 13, 28, 24, 30, 20, -37, 18, 22, 22, 0, 6, 9, 15, 3, 10, -8, -14, -5, -14, 4, 11, -9, -19, -13, 3, 21, 13, 4, 0, 2, -29, -32, -39, 9, 2, 5, -23, -34, -7, -6, -4, 7, 0, -20, -40, -49, -17, 13, 6, 27, 1, -18, -19, -8, -14, -12, -17, -29, -7, 4, 2, -19, 4, 1, -5, -13, -17, 11, -9, -33, -26, -28, -4, 17, -9, 0 },
    { 1, 6, -1, -14, -22, -38, -38, 26, -4, -30, -31, -9, 6, -7, -6, 5, -15, -13, -12, -10, 14, 17, 3, -14, -30, -20, -7, -5, -3, 34, 29, 14, 6, -4, 23, 17, 15, -1, -11, -31, -33, -2, 24, 23, 8, 9, -2, 15, 9, 14, 2, 8, 10, -5, -30, -2, 19, 31, 10, 18, 14, 2, 6, 21, 3, 13, 3, 11, -31, 36, 4, 16, 10, 0, -20, -23, 0, 29, -6, 8, 8, -5, -6, 39, 9, -4, -39, -56, -38, -48, 7, 31, 14, -3, -8, -30, 22, 42, 6, -20, -47, -37, -17, -22, 25, 46, 5, -11, -9, -15, -13, 11, 20, 15, -10, 1, 1, 1, 27, 24, -13, -23, -13, 6, 24, 24, 25, 3, 3, 4, 15, -5, 12, 3, -11, 9, 2, 26, 22, 41, -8, 8, 13, 34, 18, -4, -6, -13, -3, 15, 14, 13, 10, -3, 18, 3, 37, 31, 11, -6, 4, 0, 0, 5, -3, -2, -14, -1, 9, 7, -3, -4, -3, -2, 2, -6, -14, -14, -18, -43, -27, 25, 3, -8, -13, -6, 3, -14, -17, -17, -1, 18, -22, -14, 1, 8 },
    { 1, -7, 4, -16, -7, -4, -6, -20, 27, -32, -37, -12, -2, -1, 7, 11, 25, 28, 33, 29, 9, -6, -1, -5, -5, -3, 21, 7, -2, -4, 12, 13, 9, 5, -7, -8, -11, -8, -18, -28, -6, -19, -27, -5, -18, -17, -16, -37, -25, -11, 6, -5, -6, -16, 2, 3, -8, -7, -42, -17, -17, -13, -1, 6, -8, -7, -3, -14, -12, -31, -2, -11, -11, 7, -3, -4, 4, -18, -10, -6, -5, -25, -28, -44, -9, -30, -12, 14, 1, 18, 24, -5, -7, 12, -11, -6, -1, -4, -8, 19, 4, 17, 26, 34, 35, 23, 19, 9, -11, 9, 12, 45, -22, 8, 18, 11, 17, 29, 3, 28, 37, 21, 6, 0, 13, 40, -27, 12, 17, 3, 0, 14, 4, 29, 23, 11, 14, 17, 8, 8, 11, 19, 4, -16, -20, -8, -10, -23, -30, -12, -11, -4, 3, 15, 2, 5, -19, -20, -18, -24, -32, -43, -35, -42, -25, -16, -15, -23, -2, -27, -2, 1, -27, -20, -18, -16, -8, 6, 4, -7, 3, 17, 2, 8, 37, 13, -1, -3, 19, 27, 17, 17, 12, 4, 17, 5 },
    { -6, 0, 7, -8, -5, -2, -12, 4, -1, -9, -10, 0, 8, -1, 8, -7, 9, 8, 16, 15, -11, -29, -31, -30, -10, 4, 15, -4, 8, 8, -5, 10, 10, 29, 20, -2, -24, -11, -11, 3, 6, 27, -15, 27, -6, 11, 30, 36, 40, 52, 35, 14, -10, -28, -40, -6, 15, 10, 7, 13, 7, 17, 19, 27, 14, 4, -10, -16, -13, -7, 32, 25, 25, 18, 9, -1, 8, -5, 4, 19, 6, -3, 11, 18, 19, 19, 2, -13, -13, -23, -30, -6, 5, 10, 0, -18, -30, -14, 4, 1, -22, -12, -15, -15, -5, -8, -17, -11, 0, -15, -23, -17, -10, -4, -12, -12, -9, 9, -3, -22, -6, -19, 1, -3, -5, 6, 14, -19, -19, -5, -6, 8, -23, -20, -6, 7, 18, 23, 0, 18, 20, -32, 0, -11, -19, -23, -6, -8, 1, 6, 8, 10, 21, 13, -4, -19, -22, 18, 2, 13, 19, 8, 2, -12, -9, 12, 28, -27, 6, 2, 14, 20, 20, 23, 26, 27, 22, 12, 22, 8, 15, -14, 5, 18, 0, 11, 81, 80, 69, 79, 78, 79, 62, 39, 21, 2 },
    { 1, -4, 5, -9, 10, 5, 0, 5, -24, 22, 21, 6, -9, -5, 9, -3, 6, 4, 2, -5, -19, -4, -4, 8, 12, 35, 4, -6, 2, -23, -3, 15, 11, 4, 1, -2, 8, 6, 25, 23, 21, 19, -19, -19, 13, 10, 17, -2, -28, -22, -4, -4, -2, 15, 40, 17, -3, 6, 11, 8, 14, 2, -13, -38, -10, 3, 9, -9, 24, 11, 0, -11, -2, 6, 21, 14, 12, -11, -2, -6, -16, -9, -14, 4, 18, -2, 3, 15, 16, 24, 24, 1, 12, -4, 9, 2, 9, -25, 13, 10, -2, 15, 14, 13, 2, 9, 10, 11, -3, 2, -15, -32, -10, -8, -10, 13, 22, 0, 7, 34, 12, 3, 4, 5, 2, -24, -33, 13, 0, 2, -13, -1, 12, 13, -5, -3, 5, -1, 3, -11, -12, -17, -17, -6, -3, -4, -4, 7, -5, -7, -7, -13, -36, -24, 4, -45, -4, -17, -5, -2, 0, 10, 18, 7, -1, -16, -20, 3, 9, -35, -38, -25, -17, -3, -7, 7, -4, -4, -19, -18, -25, -10, -4, -15, -21, -25, -45, -49, -45, -57, -45, -45, -44, -10, -17, 0 },
    { 2, 7, 5, 15, 26, 6, -1, 13, 9, 48, 28, 20, -4, 8, -6, -7, 2, 30, 27, 10, 7, 6, -3, -1, -6, 18, 6, 2, 1, 15, 34, 13, 2, -9, -9, -11, -16, -9, 2, -3, -12, 3, -32, -14, 5, -22, -36, -2, -7, -6, -12, -9, -6, 0, -22, -4, -22, -10, -2, -23, -14, 14, 3, -6, -10, 0, -4, -9, -56, -27, -15, -21, 4, -13, 1, 3, -16, -4, -7, 9, 3, -17, -41, -38, -26, -26, 3, 1, 17, -10, -6, 5, -4, 0, 5, 10, 4, -11, -20, 5, 8, 16, 23, -2, 29, 22, 8, 2, 6, 2, -6, 45, 4, 1, -3, -7, -6, 8, 17, 24, -1, -9, -4, 1, 9, 29, -25, -15, -23, -16, -11, -8, 7, 13, 6, 16, 22, 12, 24, 21, -16, 13, -11, 0, 10, 7, 6, 16, 14, 24, 19, 13, 10, -2, 12, 20, 16, 3, 24, 5, -8, -14, -8, 9, 27, 11, -5, -4, -3, -37, -31, 1, -7, -19, -21, -29, -30, -21, -2, 0, 9, 21, -8, 2, 33, 27, 4, 12, 5, 5, -5, -33, -13, -33, 20, -6 },
    { -1, -5, -1, -6, -8, 3, 0, 8, -10, 38, 35, 16, -5, -5, 1, 12, 10, -12, 13, -9, -28, -28, -5, 19, 13, 14, 9, 25, 4, 14, 25, 12, -9, -21, -26, -25, -35, -27, -16, 0, -2, -9, -10, 27, -7, -3, -3, -1, -2, -5, 2, -5, 0, 3, -2, 0, 24, 13, -13, -12, -4, -21, 5, 26, 34, 32, 28, 16, 11, -2, 24, 25, -23, -13, -23, -24, 15, 32, 21, 15, 14, 13, 34, 17, 9, 32, -31, -5, -9, 7, 10, 10, -14, -29, -47, -77, -21, 23, 18, 13, 12, 3, 3, 12, 2, -3, -2, -1, -5, -64, -47, -22, -14, -13, 24, 20, -2, -2, 1, 2, 10, 11, -15, -70, -27, -11, 25, -35, 7, 15, -1, 12, 31, 8, 2, -1, -40, -41, -22, 24, -4, -38, -28, -5, 2, -2, 19, -1, -23, -21, -52, -27, -8, -5, 3, -20, -1, -1, -3, 3, -10, -19, -26, -43, -21, -6, -23, 23, 8, 5, 43, -1, 7, -8, -1, -15, -19, -28, -32, -6, 19, 6, 2, 2, -8, -13, 20, 23, 27, 23, 14, -4, -7, 5, 0, 0 },
    { -8, 4, -9, -9, -3, -6, -7, -15, -12, -5, -11, -1, -1, -5, -3, 5, 22, -4, 11, -2, -4, -10, -6, 9, 19, 5, 9, -10, 3, -7, 8, 14, 4, 27, 19, 14, 20, 21, 8, 11, 5, 14, 12, -9, 3, -4, 7, -4, 13, 10, 9, 0, 3, -2, 8, 14, -19, -3, -5, -5, 10, 11, -1, -10, -6, -8, -8, -4, -4, 11, -24, 3, -8, 4, 1, 0, 5, 7, 10, 1, -8, -26, -31, 4, -18, -33, -16, -10, -6, 7, 41, 45, 24, 13, -7, -20, -23, 10, 19, -16, -50, -44, -34, 6, 23, 6, -3, -3, -3, 22, 15, -14, 13, 18, -18, -58, -101, -90, -57, -21, -8, 7, 13, 12, 10, -45, -12, 46, 26, 5, -12, -37, -44, -12, -6, 2, 17, -8, -19, -46, 8, 8, 19, 26, 31, 31, 8, 0, -8, -9, -1, -17, -36, -19, -12, 16, 19, 7, 10, 16, 12, 0, 1, -11, -18, -20, -25, -2, 4, 31, 35, 36, 20, 11, -1, -11, 12, -25, -17, 0, -19, -7, 6, 11, 33, 19, 34, 25, 20, 36, 26, 24, 21, 7, 10, -2 },
    { 9, -2, 0, -12, 16, 0, 5, -4, -14, 13, 14, -12, -5, -3, 5, -7, 16, 15, -12, 5, -8, 4, -4, 16, 31, 58, -6, 11, -2, -12, -15, -3, -1, 6, 2, -7, -19, -3, 8, 29, 56, 27, -12, -40, -6, -8, 9, 3, 1, 3, -1, -3, 3, 10, 41, 68, -25, -18, -4, 7, 7, -11, -36, -30, -9, -2, 3, 3, 46, 17, -36, -36, 1, 15, 40, 17, -24, -33, -10, -12, -21, -10, 17, -2, -6, -26, -1, 27, 33, 25, 3, -4, 8, 7, 5, 13, -15, -36, 9, -10, 7, 10, 32, 23, 4, -2, 20, 6, -8, 1, -25, -31, -13, -25, -32, 5, 18, 19, 19, -5, 18, 11, -2, -15, -12, -25, -29, -28, -21, -11, 10, 11, 35, -1, 0, 5, -4, -17, -5, -37, 0, -28, -23, -31, -16, -2, 7, 4, -1, 2, 1, 7, -10, -28, -4, -30, -39, -33, -17, -12, -7, 13, 8, 12, 16, 0, 5, 2, -1, -8, -16, -15, -5, 3, -7, 9, 5, 19, 11, 17, -25, -10, -5, -4, -11, -10, 2, -2, 0, -7, -22, -19, -29, -38, -21, 7 },
    { -8, 4, -3, 12, 10, 7, 23, 20, 32, 17, -7, 1, 0, 6, -5, 11, 12, 3, 3, -11, -1, -4, 11, 26, 15, -5, 4, 16, 9, -6, 10, -12, 1, -1, -2, 3, 1, 8, 8, 10, 5, 6, 19, -10, -7, 3, 1, 10, 5, 10, -8, 13, 22, 31, 31, 29, -10, -25, -28, -5, -2, 19, 20, -5, -15, -12, -4, 13, 27, 21, -33, -1, -10, 2, 0, 6, 17, 0, -22, -34, -57, -79, -18, 33, -18, -5, -6, 1, -7, -11, 15, 4, -2, -6, -33, -78, -94, 18, 9, -21, -27, -8, 12, 3, 10, 3, -4, -3, -5, -13, -27, -19, 20, 23, -15, -19, -9, 2, 3, -9, -17, 11, 9, -1, 3, -7, -6, 41, -6, -19, -36, -47, -31, -6, 4, 14, 23, 7, 8, -29, -9, 9, 13, -7, 15, 7, 7, 9, 12, 34, 31, 42, 34, -5, -1, 18, 38, 10, 8, 5, 8, 13, 13, 20, 15, 17, -5, 17, -6, 22, 16, 27, 25, 22, 13, 5, 16, 3, 15, 26, 13, 21, -7, 7, 0, -8, -4, 1, -2, 17, 33, -3, 16, 12, 6, -3 },
    { -6, 2, 7, 18, 23, 32, 24, 2, 51, 39, 18, 16, 0, 4, -2, -2, -4, 9, 21, 34, 22, 16, 25, 39, 20, 34, 36, 24, -11, -12, -43, -28, -11, 18, 15, 12, 39, 28, 14, 16, 17, 48, -27, -11, -22, -4, 7, 8, 14, 31, 24, 15, 10, 18, 17, 2, -5, -24, -14, 3, 12, 16, -1, -10, -16, -17, -15, -2, 6, -8, -25, -39, -2, 15, 5, 3, -13, -43, -38, -28, -33, -29, 33, -2, -26, 4, -21, -12, -4, 12, 3, -26, -16, -8, -12, -3, 7, 1, -1, -11, -29, -8, -5, 6, 9, -3, -16, -9, -4, -1, 34, 32, -23, 3, -10, -6, -23, 12, 19, -18, -11, -22, 3, -5, 25, 19, -25, -12, 11, 10, -4, -1, -7, -13, 9, 4, -13, -4, 15, 1, -4, 12, 5, 4, 24, 23, 29, 29, 19, 6, 8, 29, 18, 11, -23, 12, -8, 4, 22, 26, 36, 29, 18, 10, 15, 34, 23, -10, -1, -15, -18, -8, 10, 11, 13, 19, 20, 31, 19, 29, 31, -9, -5, 0, -8, -21, -34, 6, 9, -24, -2, -10, 3, -11, 10, 2 },
    { 8, 2, -2, -27, -16, -33, -39, -24, 2, -33, -37, -29, 1, 2, 2, -7, 1, 9, 12, 29, 12, 6, -13, -20, -15, -6, 5, 3, 2, 11, -6, 8, 13, 8, 0, 3, 8, -1, 12, 36, 25, -3, 19, 0, 22, 10, 3, -11, -6, -11, -35, -31, -12, 14, 39, 21, 3, 12, 7, -9, -6, -8, 1, -9, -4, 1, 19, 9, 3, -2, -4, 4, -8, -5, -25, -25, -4, -26, 8, 2, -5, -5, -12, -29, 2, -12, -21, -7, -19, 18, 27, -20, -8, -11, -1, -17, 20, 1, 15, 17, 8, 11, 9, 12, 20, 13, 4, -3, -10, -8, 6, 52, 8, 37, 5, 16, 3, 4, 19, 16, 14, 2, 6, 12, 11, 31, -25, 31, 18, 8, -3, 1, 16, 18, 27, 1, 12, 0, -7, 11, 5, 39, 15, -5, 11, 14, 14, 9, 14, 8, 13, 12, -11, 21, -12, 27, -9, -10, 6, 18, 11, -3, 6, 12, 16, 7, -13, -11, 6, -15, -31, -46, -33, -30, -22, -3, -16, -11, -16, -10, 14, -2, -1, -1, -14, -50, -69, -69, -77, -74, -43, -51, -57, -35, -6, 1 },
    { -8, 5, 8, 21, 11, 9, -1, 6, 3, 42, 37, 16, -2, 9, 3, -3, 0, 27, -1, 6, 12, 27, 12, 12, 25, 21, 4, 3, 6, -15, 0, 3, 11, -10, -9, -7, -13, -14, -10, -5, -30, -35, -25, 12, 0, 17, 2, -13, 1, -1, -1, -17, -17, -14, -35, -3, 32, 9, 13, 8, -2, 1, 1, 2, -15, -27, -27, -3, -13, -8, 23, 15, -5, -3, -7, 11, 19, 16, 11, -2, -15, -12, -29, -26, 24, 13, -4, 3, 3, 30, 2, 16, 35, 16, 2, -10, -26, -17, 11, 16, -8, 0, 4, 29, 0, 5, 32, 27, 14, 22, -35, -15, -9, -15, 5, 1, -2, 7, -21, 17, 32, 14, 15, -2, 0, 4, 10, -4, -5, -28, -27, -26, -10, 16, -12, -18, -29, -31, 8, 23, -14, -18, -19, -33, -28, -10, 4, -9, -21, -38, -57, -42, -11, -7, 1, -49, -44, -11, 6, 1, -13, -20, -8, -20, -17, -35, -16, -12, -7, -17, -25, -2, 4, 3, -10, 3, 8, 11, 17, 3, -11, -3, 9, 7, -8, 22, 39, 14, 9, 31, 10, 22, 6, 11, 5, 9 }
    };
    
    wire dense1_en = enable;
    reg dense1_done = 0;

    
    dense_layer #(.NEURON_NB(32),.IN_SIZE(196), .WIDTH(8)) dense_layer1(.clk(clk), .layer_en(dense1_en), .reset(reset),
                                                                        .in_data(pooled_img), .weights(W_ARRAY_L2), .biases(B_ARRAY_L2),
                                                                        .neuron_out(dense1_res), .layer_done(dense1_done)); //Dense layer
    
    relu relu_activation[31:0] (.data_in(dense1_res), .data_out(relu_res)); //ReLu activation
    
    assign layer_out = relu_res;               
    assign layer_done = dense1_done;

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.12.2022 09:16:01
// Design Name: 
// Module Name: dense_layer2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/**********
* 1st dense layer implementation (output layer)
*
* Inputs: clk => clock signal, enable => enable signal, 
*         reset => active high sync reset, in_data => in vector, 
*
* Outputs: layer_out => dense layer output
*          layer_done => done signal
* 
***********/

module dense_layer2(
    input clk,
    input enable,
    input reset,
    input signed [15:0] in_data [0:31],
    output signed [15:0] layer_out [0:9],
    output layer_done
    );
    
    reg signed [31:0] dense2_res [0:9];
    reg signed [15:0] relu_res [0:9];
  
    //Biases and weights
    localparam signed [7:0] B_ARRAY_L3 [0:9] = '{ -11, 10, 14, -23, -1, 8, 0, 13, 1, -11 };
    
    localparam signed [7:0] W_ARRAY_L3 [0:9] [0:31] = '{
    { 33, -57, -6, -23, -11, -48, -53, 46, -54, -24, 4, 9, -2, -40, -29, 20, -6, 45, -85, 2, -57, 45, 40, -21, -23, -2, -105, -19, -40, 28, -7, 15 },
    { 30, 34, 29, -19, -12, -47, 50, -69, 64, -25, 38, 35, -43, 19, -17, -61, 62, -31, -30, -69, 43, -67, -60, 5, 46, -1, -50, -64, 39, -39, -28, -28 },
    { 2, -48, 30, 33, 69, -11, 28, -1, 28, 25, -22, 58, -11, -120, -6, -28, -72, -12, -33, -4, 1, 81, 21, -22, 24, -100, -59, -59, -20, 27, 37, 39 },
    { -37, 61, -6, -19, -5, 60, 14, 8, 28, -29, -106, 53, 32, -18, -27, -16, -1, -45, 43, 40, 18, -28, 25, -37, -7, -23, 52, -45, 16, -28, 6, -53 },
    { -9, 57, 20, 19, -96, -25, -47, 19, 43, -19, 8, -68, -37, 37, 28, -8, 13, -15, 17, -40, -33, 2, -100, 35, 5, -52, 12, 34, -75, -92, 30, 17 },
    { 16, -8, -127, -69, 28, -82, 29, -47, -7, -19, -11, -55, -10, 37, -46, -14, 26, -1, 39, 35, -37, -5, 10, -20, -35, 84, 55, 13, 37, 25, -5, -36 },
    { 40, 29, -74, -1, -16, 71, -91, -13, -92, 24, 32, -15, -5, -12, -73, -70, 0, -25, -85, 38, -63, 2, -53, 36, 39, 4, -93, 24, 26, 19, 12, 37 },
    { -40, -42, -10, 45, 26, 8, 25, 8, -33, -40, -32, 34, -40, -38, 32, 19, 42, -20, -18, 41, 21, -41, 24, 7, -25, 37, -93, -32, -56, -52, -48, 55 },
    { 4, -73, 17, -34, 17, 0, -34, -9, -50, 10, 29, -75, 37, 10, -19, 0, -63, -1, 12, 2, 9, -63, 7, 40, -12, -54, -17, 26, -10, -5, -7, -89 },
    { -82, -31, 23, -61, -34, 18, -52, -24, -1, 12, 29, -74, -11, 14, 34, 33, 23, -13, -21, -98, -48, 32, 26, -35, 7, 3, 68, 14, -25, -11, -86, 27 }
    };
    
    wire dense2_en = enable;
    reg dense2_done = 0;

    
  dense_layer #(.NEURON_NB(10),.IN_SIZE(32), .WIDTH(8)) dense_layer2(.clk(clk), .layer_en(dense2_en), .reset(reset),
                                                                     .in_data(in_data), .weights(W_ARRAY_L3), .biases(B_ARRAY_L3),
                                                                     .neuron_out(dense2_res), .layer_done(dense2_done)); //Dense layer

    relu relu_activation[9:0] (.data_in(dense2_res), .data_out(relu_res)); //ReLu activation
    
    assign layer_out = relu_res;               
    assign layer_done = dense2_done;

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.12.2022 10:34:30
// Design Name: 
// Module Name: neural_network
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/**********
* Neural Network implementation
*
* Inputs: clk => clock signal, enable => NN enable signal, img => in vector, 
*
* Outputs: digit out => handwritten digit
*          NN_done => done signal
* 
***********/

module neural_network(
    input clk,
    input enable,
    input reset,
    input [7:0] img [0:783],
    output [7:0] digit_out,
    output NN_done
    );
    
    /* Average pooling layer */
    
    reg pool_enable;
    wire finished_pool;
    reg signed [15:0] pool [0:195];
    
    // Pixel value registers
    wire signed [7:0] pool_in1;
    wire signed [7:0] pool_in2;
    wire signed [7:0] pool_in3;
    wire signed [7:0] pool_in4;
    wire signed [7:0] pool_final;
    
    // Pixel address registers
    reg [15:0] pool_in1_addr;
    reg [15:0] pool_in2_addr;
    reg [15:0] pool_in3_addr;
    reg [15:0] pool_in4_addr;
    reg [15:0] pool_final_addr = 0;
    reg [15:0] pool_addr = 0;
    reg [15:0] pool_row = 0;
    
    // Initialize addresses
    initial
    begin
        pool_in1_addr <= 8'b0000_0000;
        pool_in2_addr <= 8'b0000_0001;
        pool_in3_addr <= 8'b0001_1100;
        pool_in4_addr <= 8'b0001_1101;
        pool_enable <= 1'b1;
    end
    
    avg_pooling AvgPooling(clk,pool_enable,pool_in1,pool_in2,pool_in3,pool_in4,pool_final,finished_pool);
    
    // Load pixel values
    assign pool_in1 = ((img[pool_in1_addr]));
    assign pool_in2 = ((img[pool_in2_addr]));
    assign pool_in3 = ((img[pool_in3_addr]));
    assign pool_in4 = ((img[pool_in4_addr]));
    
    always @(posedge clk) begin
    if(reset) begin
        pool_in1_addr <= 8'b0000_0000;
        pool_in2_addr <= 8'b0000_0001;
        pool_in3_addr <= 8'b0001_1100;
        pool_in4_addr <= 8'b0001_1101;
        pool_final_addr <= 0;
        pool_row <= 0;
        pool_addr <= 0;
        pool_enable <= 1'b1; 
    end
    else if(enable) begin
        if(finished_pool) begin // Average done
            pool[pool_final_addr] = pool_final;
            pool_addr <= pool_addr + 2; // Increment address
            pool_row <= pool_row + 2;
            if(pool_row == 28) begin // End of row, go down by 2 rows
                pool_addr <= pool_addr + pool_row;
                pool_row <= 0;
            end
            if(pool_in4_addr == 783) begin // Global averaging done
                pool_enable <= 0;
            end
            else if(pool_in4_addr != 783) begin // Update addresses
                pool_in1_addr <= pool_addr;
                pool_in2_addr <= pool_addr + 1;
                pool_in3_addr <= pool_addr + 28;
                pool_in4_addr <= pool_addr + 29;
                pool_final_addr <= pool_final_addr + 1;
            end
        end
    end       
    end
    
    /* Hidden layer */
    
    reg dense1_enable;
    wire finished_dense1;
    reg signed [15:0] dense1_res [0:31];
    initial dense1_enable <= 0;
    
    dense_layer1 layer2 (.clk(clk), .enable(dense1_enable), .reset(reset), .pooled_img(pool), .layer_out(dense1_res), .layer_done(finished_dense1));

    always @(posedge clk) begin
        if(reset) begin
            dense1_enable <= 0;
        end
        else if(enable) begin
            if(pool_enable == 0 && finished_dense1 == 0) begin // Pooling done
                dense1_enable <= 1;
            end
            else dense1_enable <= 0; // Hidden layer done
        end
    end
    
    /* Output layer */
    
    reg dense2_enable;
    wire finished_dense2;
    reg signed [15:0] dense2_res [0:9];
    initial dense2_enable <= 0;

    dense_layer2 layer3 (.clk(clk), .enable(dense2_enable), .reset(reset), .in_data(dense1_res), .layer_out(dense2_res), .layer_done(finished_dense2));

    always @(posedge clk) begin
        if(reset) begin
            dense2_enable <= 0;
        end
        else if(enable) begin
            if(pool_enable == 0 && finished_dense1 == 1 && finished_dense2 == 0) begin // Previous layers done
                dense2_enable <= 1;
            end
            else dense2_enable <= 0; // Output layer done
        end
    end
    
    /* Handwritten digit selection layer */
    
    reg max_enable;
    wire digit_recog_done;
    reg [7:0] digit;
    
    initial max_enable <= 0;
    
    select_max last_layer (.clk(clk), .enable(max_enable), .reset(reset), .in_data(dense2_res), .digit(digit), .layer_done(digit_recog_done));
        
    always @(posedge clk) begin
        if(reset) begin
            max_enable <= 0;
        end
        else if(enable) begin
            if(finished_dense2 == 1) begin // Output layer done
                max_enable <= 1;
            end
            else max_enable <= 0;
        end
    end
    
    assign digit_out = digit;
    assign NN_done = digit_recog_done;
    
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.12.2022 23:18:14
// Design Name: 
// Module Name: neuron
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


/**********
* Single neuron implementation
*
* Parameters: IN_SIZE => The input vector size
*             WIDTH => The width of the weights and biases
*
* Inputs: clk => clock signal, en => enable signal,
*         in_data => in vector, reset => active high sync reset
*         weights => neuron weights, bias => neuron bias
*
* Outputs: neuron_out => neuron value after activation
*          neuron_done => done signal
* 
***********/


module neuron #(parameter IN_SIZE=196, WIDTH = 8)(
    input clk,
    input en,
    input reset,
    input signed [2*WIDTH-1:0] in_data[0:IN_SIZE-1],
    input signed[WIDTH-1:0] weight[0:IN_SIZE-1],
    input signed[WIDTH-1:0] bias,
    output signed[4*WIDTH-1:0] neuron_out,
    output neuron_done
    );
    
    integer addr = 0;
    reg done = 0;
    
    reg signed [4*WIDTH-1:0] product = 0;
    reg signed [4*WIDTH-1:0] out = 0;
    
    always @(posedge clk) begin
        if(reset) begin 
            done <= 0;
            addr <= 0;
        end
        else if(en) begin
            if(addr < IN_SIZE-1) begin
                product <= in_data[addr]*weight[addr]; //Calculate weighted input
                out <= out+product; //Sum each weighted input
               
            end
            if(addr == IN_SIZE-1) begin //Neuron output available
                done <= 1;
            end else begin
                addr <= addr + 1'b1;
                done <= 0;
            end
        end
    end
    
    assign neuron_out = out + bias; //Add bias
    assign neuron_done = done;
    
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.01.2023 15:38:43
// Design Name: 
// Module Name: relu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


/**********
* Relu activation function implementation
*
* Parameters: WIDTH => The width used in the NN
*
* Inputs: data_in => in element, 
*
* Outputs: data_out => relu output (ie data_in if >0, else 0)
* 
***********/


module relu #(parameter WIDTH = 8)(
    input signed [4*WIDTH-1:0] data_in,
    output signed [2*WIDTH-1:0] data_out
    );
    
    wire signed [4*WIDTH-1:0] temp;
    
    assign temp = (data_in > 0)? data_in:0; //Take data_in if > 0, 0 else
    assign data_out = temp >> 8; //Rescale element and store into data_out
    
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.01.2023 22:59:45
// Design Name: 
// Module Name: select_max
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/**********
* Module to select the maximum between last layer outputs
*
* Inputs: clk => clock signal, enable => enable signal,
*         reset => active high sync reset, in_data => input array, 
*
* Outputs: digit => Index of max element (ie handwritten digit)
*          layer_done => done signal
* 
***********/

module select_max # (parameter NEURON_NB=10, WIDTH=8)(
    input clk,
    input enable,
    input reset,
    input signed[2*WIDTH-1:0] in_data [0:NEURON_NB-1],
    output [WIDTH-1:0] digit,
    output layer_done
    );
    
    integer i = 0;
    reg signed [2*WIDTH-1:0] max = 0;
    reg signed [WIDTH-1:0] index = 0;
    reg done = 0;
    
    always @(posedge clk) begin
        if(reset) begin
            done <= 0;
            i <= 0;
            max <= 0;
            index <= 0;
        end
        else if(enable) begin
            if (in_data[i] >= max) begin //Update maximum and max index
                    max <= in_data[i]; 
                    index <= i;
                end
            if(i < 10) i <= i + 1;
                else done <= 1;
        end
    end
    
    assign digit = index;
    assign layer_done = done;
    
endmodule

